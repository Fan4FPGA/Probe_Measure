library verilog;
use verilog.vl_types.all;
entity altmult_accum is
    generic(
        width_a         : integer := 2;
        width_b         : integer := 2;
        width_result    : integer := 5;
        input_reg_a     : string  := "CLOCK0";
        input_aclr_a    : string  := "ACLR3";
        input_reg_b     : string  := "CLOCK0";
        input_aclr_b    : string  := "ACLR3";
        port_addnsub    : string  := "PORT_CONNECTIVITY";
        addnsub_reg     : string  := "CLOCK0";
        addnsub_aclr    : string  := "ACLR3";
        addnsub_pipeline_reg: string  := "CLOCK0";
        addnsub_pipeline_aclr: string  := "ACLR3";
        accum_direction : string  := "ADD";
        accum_sload_reg : string  := "CLOCK0";
        accum_sload_aclr: string  := "ACLR3";
        accum_sload_pipeline_reg: string  := "CLOCK0";
        accum_sload_pipeline_aclr: string  := "ACLR3";
        representation_a: string  := "UNSIGNED";
        port_signa      : string  := "PORT_CONNECTIVITY";
        sign_reg_a      : string  := "CLOCK0";
        sign_aclr_a     : string  := "ACLR3";
        sign_pipeline_reg_a: string  := "CLOCK0";
        sign_pipeline_aclr_a: string  := "ACLR3";
        port_signb      : string  := "PORT_CONNECTIVITY";
        representation_b: string  := "UNSIGNED";
        sign_reg_b      : string  := "CLOCK0";
        sign_aclr_b     : string  := "ACLR3";
        sign_pipeline_reg_b: string  := "CLOCK0";
        sign_pipeline_aclr_b: string  := "ACLR3";
        multiplier_reg  : string  := "CLOCK0";
        multiplier_aclr : string  := "ACLR3";
        output_reg      : string  := "CLOCK0";
        output_aclr     : string  := "ACLR3";
        lpm_type        : string  := "altmult_accum";
        lpm_hint        : string  := "UNUSED";
        extra_multiplier_latency: integer := 0;
        extra_accumulator_latency: integer := 0;
        dedicated_multiplier_circuitry: string  := "AUTO";
        dsp_block_balancing: string  := "AUTO";
        intended_device_family: string  := "Stratix";
        accum_round_aclr: string  := "ACLR3";
        accum_round_pipeline_aclr: string  := "ACLR3";
        accum_round_pipeline_reg: string  := "CLOCK0";
        accum_round_reg : string  := "CLOCK0";
        accum_saturation_aclr: string  := "ACLR3";
        accum_saturation_pipeline_aclr: string  := "ACLR3";
        accum_saturation_pipeline_reg: string  := "CLOCK0";
        accum_saturation_reg: string  := "CLOCK0";
        accum_sload_upper_data_aclr: string  := "ACLR3";
        accum_sload_upper_data_pipeline_aclr: string  := "ACLR3";
        accum_sload_upper_data_pipeline_reg: string  := "CLOCK0";
        accum_sload_upper_data_reg: string  := "CLOCK0";
        mult_round_aclr : string  := "ACLR3";
        mult_round_reg  : string  := "CLOCK0";
        mult_saturation_aclr: string  := "ACLR3";
        mult_saturation_reg: string  := "CLOCK0";
        input_source_a  : string  := "DATAA";
        input_source_b  : string  := "DATAB";
        width_upper_data: integer := 1;
        multiplier_rounding: string  := "NO";
        multiplier_saturation: string  := "NO";
        accumulator_rounding: string  := "NO";
        accumulator_saturation: string  := "NO";
        port_mult_is_saturated: string  := "UNUSED";
        port_accum_is_saturated: string  := "UNUSED";
        int_width_a     : vl_notype;
        int_width_b     : vl_notype;
        int_width_result: vl_notype;
        int_extra_width : vl_notype;
        diff_width_a    : vl_notype;
        diff_width_b    : vl_notype;
        sat_for_ini     : vl_notype;
        mult_round_for_ini: vl_notype;
        bits_to_round   : vl_notype;
        sload_for_limit : vl_notype;
        accum_sat_for_limit: vl_notype
    );
    port(
        dataa           : in     vl_logic_vector;
        datab           : in     vl_logic_vector;
        scanina         : in     vl_logic_vector;
        scaninb         : in     vl_logic_vector;
        sourcea         : in     vl_logic;
        sourceb         : in     vl_logic;
        accum_sload_upper_data: in     vl_logic_vector;
        addnsub         : in     vl_logic;
        accum_sload     : in     vl_logic;
        signa           : in     vl_logic;
        signb           : in     vl_logic;
        clock0          : in     vl_logic;
        clock1          : in     vl_logic;
        clock2          : in     vl_logic;
        clock3          : in     vl_logic;
        ena0            : in     vl_logic;
        ena1            : in     vl_logic;
        ena2            : in     vl_logic;
        ena3            : in     vl_logic;
        aclr0           : in     vl_logic;
        aclr1           : in     vl_logic;
        aclr2           : in     vl_logic;
        aclr3           : in     vl_logic;
        result          : out    vl_logic_vector;
        overflow        : out    vl_logic;
        scanouta        : out    vl_logic_vector;
        scanoutb        : out    vl_logic_vector;
        mult_round      : in     vl_logic;
        mult_saturation : in     vl_logic;
        accum_round     : in     vl_logic;
        accum_saturation: in     vl_logic;
        mult_is_saturated: out    vl_logic;
        accum_is_saturated: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width_a : constant is 1;
    attribute mti_svvh_generic_type of width_b : constant is 1;
    attribute mti_svvh_generic_type of width_result : constant is 1;
    attribute mti_svvh_generic_type of input_reg_a : constant is 1;
    attribute mti_svvh_generic_type of input_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of input_reg_b : constant is 1;
    attribute mti_svvh_generic_type of input_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of port_addnsub : constant is 1;
    attribute mti_svvh_generic_type of addnsub_reg : constant is 1;
    attribute mti_svvh_generic_type of addnsub_aclr : constant is 1;
    attribute mti_svvh_generic_type of addnsub_pipeline_reg : constant is 1;
    attribute mti_svvh_generic_type of addnsub_pipeline_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_direction : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_reg : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_pipeline_reg : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_pipeline_aclr : constant is 1;
    attribute mti_svvh_generic_type of representation_a : constant is 1;
    attribute mti_svvh_generic_type of port_signa : constant is 1;
    attribute mti_svvh_generic_type of sign_reg_a : constant is 1;
    attribute mti_svvh_generic_type of sign_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of sign_pipeline_reg_a : constant is 1;
    attribute mti_svvh_generic_type of sign_pipeline_aclr_a : constant is 1;
    attribute mti_svvh_generic_type of port_signb : constant is 1;
    attribute mti_svvh_generic_type of representation_b : constant is 1;
    attribute mti_svvh_generic_type of sign_reg_b : constant is 1;
    attribute mti_svvh_generic_type of sign_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of sign_pipeline_reg_b : constant is 1;
    attribute mti_svvh_generic_type of sign_pipeline_aclr_b : constant is 1;
    attribute mti_svvh_generic_type of multiplier_reg : constant is 1;
    attribute mti_svvh_generic_type of multiplier_aclr : constant is 1;
    attribute mti_svvh_generic_type of output_reg : constant is 1;
    attribute mti_svvh_generic_type of output_aclr : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of lpm_hint : constant is 1;
    attribute mti_svvh_generic_type of extra_multiplier_latency : constant is 1;
    attribute mti_svvh_generic_type of extra_accumulator_latency : constant is 1;
    attribute mti_svvh_generic_type of dedicated_multiplier_circuitry : constant is 1;
    attribute mti_svvh_generic_type of dsp_block_balancing : constant is 1;
    attribute mti_svvh_generic_type of intended_device_family : constant is 1;
    attribute mti_svvh_generic_type of accum_round_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_round_pipeline_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_round_pipeline_reg : constant is 1;
    attribute mti_svvh_generic_type of accum_round_reg : constant is 1;
    attribute mti_svvh_generic_type of accum_saturation_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_saturation_pipeline_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_saturation_pipeline_reg : constant is 1;
    attribute mti_svvh_generic_type of accum_saturation_reg : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_upper_data_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_upper_data_pipeline_aclr : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_upper_data_pipeline_reg : constant is 1;
    attribute mti_svvh_generic_type of accum_sload_upper_data_reg : constant is 1;
    attribute mti_svvh_generic_type of mult_round_aclr : constant is 1;
    attribute mti_svvh_generic_type of mult_round_reg : constant is 1;
    attribute mti_svvh_generic_type of mult_saturation_aclr : constant is 1;
    attribute mti_svvh_generic_type of mult_saturation_reg : constant is 1;
    attribute mti_svvh_generic_type of input_source_a : constant is 1;
    attribute mti_svvh_generic_type of input_source_b : constant is 1;
    attribute mti_svvh_generic_type of width_upper_data : constant is 1;
    attribute mti_svvh_generic_type of multiplier_rounding : constant is 1;
    attribute mti_svvh_generic_type of multiplier_saturation : constant is 1;
    attribute mti_svvh_generic_type of accumulator_rounding : constant is 1;
    attribute mti_svvh_generic_type of accumulator_saturation : constant is 1;
    attribute mti_svvh_generic_type of port_mult_is_saturated : constant is 1;
    attribute mti_svvh_generic_type of port_accum_is_saturated : constant is 1;
    attribute mti_svvh_generic_type of int_width_a : constant is 3;
    attribute mti_svvh_generic_type of int_width_b : constant is 3;
    attribute mti_svvh_generic_type of int_width_result : constant is 3;
    attribute mti_svvh_generic_type of int_extra_width : constant is 3;
    attribute mti_svvh_generic_type of diff_width_a : constant is 3;
    attribute mti_svvh_generic_type of diff_width_b : constant is 3;
    attribute mti_svvh_generic_type of sat_for_ini : constant is 3;
    attribute mti_svvh_generic_type of mult_round_for_ini : constant is 3;
    attribute mti_svvh_generic_type of bits_to_round : constant is 3;
    attribute mti_svvh_generic_type of sload_for_limit : constant is 3;
    attribute mti_svvh_generic_type of accum_sat_for_limit : constant is 3;
end altmult_accum;
