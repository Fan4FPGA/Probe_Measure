library verilog;
use verilog.vl_types.all;
entity cycloneiii_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end cycloneiii_routing_wire;
